/*
 Copyright 2013 Ray Salemi

 Licensed under the Apache License, Version 2.0 (the "License");
 you may not use this file except in compliance with the License.
 You may obtain a copy of the License at

 http://www.apache.org/licenses/LICENSE-2.0

 Unless required by applicable law or agreed to in writing, software
 distributed under the License is distributed on an "AS IS" BASIS,
 WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 See the License for the specific language governing permissions and
 limitations under the License.
 */
class add_sequence_item extends sequence_item;
   `uvm_object_utils(add_sequence_item)

   function new(input string name = "add_sequence_item");
      super.new(name);
   endfunction

   constraint add_only {op == add_op;}

endclass : add_sequence_item
